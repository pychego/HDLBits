// 驱动74hc595芯片
// 功能： 将并行16位数据（sel和seg）转化为串行数据

module HC95driver (
    input clk,
    input reset_n,
    input[15:0] data,
    output 
);
    
endmodule